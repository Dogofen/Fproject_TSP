-- nios2_c.vhd

-- Generated using ACDS version 13.1 162 at 2014.06.22.14:25:00

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity nios2_c is
	port (
		clk_clk                           : in  std_logic                     := '0';             --                        clk.clk
		reset_reset_n                     : in  std_logic                     := '0';             --                      reset.reset_n
		key_external_connection_export    : in  std_logic_vector(3 downto 0)  := (others => '0'); --    key_external_connection.export
		ledg_external_connection_export   : out std_logic_vector(7 downto 0);                     --   ledg_external_connection.export
		to_hex_external_connection_export : out std_logic_vector(13 downto 0)                     -- to_hex_external_connection.export
	);
end entity nios2_c;

architecture rtl of nios2_c is
	component nios2_c_cpu is
		port (
			clk                                   : in  std_logic                     := 'X';             -- clk
			reset_n                               : in  std_logic                     := 'X';             -- reset_n
			reset_req                             : in  std_logic                     := 'X';             -- reset_req
			d_address                             : out std_logic_vector(24 downto 0);                    -- address
			d_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                                : out std_logic;                                        -- read
			d_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_write                               : out std_logic;                                        -- write
			d_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			d_burstcount                          : out std_logic_vector(3 downto 0);                     -- burstcount
			d_readdatavalid                       : in  std_logic                     := 'X';             -- readdatavalid
			jtag_debug_module_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                             : out std_logic_vector(18 downto 0);                    -- address
			i_read                                : out std_logic;                                        -- read
			i_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			i_burstcount                          : out std_logic_vector(3 downto 0);                     -- burstcount
			i_readdatavalid                       : in  std_logic                     := 'X';             -- readdatavalid
			dcm0_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			dcm0_waitrequest                      : in  std_logic                     := 'X';             -- waitrequest
			dcm0_readdatavalid                    : in  std_logic                     := 'X';             -- readdatavalid
			dcm0_address                          : out std_logic_vector(18 downto 0);                    -- address
			dcm0_read                             : out std_logic;                                        -- read
			dcm0_clken                            : out std_logic;                                        -- clken
			dcm0_write                            : out std_logic;                                        -- write
			dcm0_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			dcm0_byteenable                       : out std_logic_vector(3 downto 0);                     -- byteenable
			icm0_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			icm0_waitrequest                      : in  std_logic                     := 'X';             -- waitrequest
			icm0_readdatavalid                    : in  std_logic                     := 'X';             -- readdatavalid
			icm0_address                          : out std_logic_vector(16 downto 0);                    -- address
			icm0_read                             : out std_logic;                                        -- read
			icm0_clken                            : out std_logic;                                        -- clken
			d_irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			jtag_debug_module_resetrequest        : out std_logic;                                        -- reset
			jtag_debug_module_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			jtag_debug_module_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_debug_module_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			jtag_debug_module_read                : in  std_logic                     := 'X';             -- read
			jtag_debug_module_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_debug_module_waitrequest         : out std_logic;                                        -- waitrequest
			jtag_debug_module_write               : in  std_logic                     := 'X';             -- write
			jtag_debug_module_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			no_ci_readra                          : out std_logic                                         -- readra
		);
	end component nios2_c_cpu;

	component nios2_c_tightly_coupled_instruction_memory is
		port (
			clk         : in  std_logic                     := 'X';             -- clk
			address     : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			clken       : in  std_logic                     := 'X';             -- clken
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset       : in  std_logic                     := 'X';             -- reset
			reset_req   : in  std_logic                     := 'X';             -- reset_req
			address2    : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			chipselect2 : in  std_logic                     := 'X';             -- chipselect
			clken2      : in  std_logic                     := 'X';             -- clken
			write2      : in  std_logic                     := 'X';             -- write
			readdata2   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata2  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable2 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			clk2        : in  std_logic                     := 'X';             -- clk
			reset2      : in  std_logic                     := 'X';             -- reset
			reset_req2  : in  std_logic                     := 'X'              -- reset_req
		);
	end component nios2_c_tightly_coupled_instruction_memory;

	component nios2_c_pll_100 is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component nios2_c_pll_100;

	component nios2_c_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component nios2_c_jtag_uart;

	component nios2_c_sysid_qsys_0 is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component nios2_c_sysid_qsys_0;

	component altera_avalon_mm_clock_crossing_bridge is
		generic (
			DATA_WIDTH          : integer := 32;
			SYMBOL_WIDTH        : integer := 8;
			ADDRESS_WIDTH       : integer := 10;
			BURSTCOUNT_WIDTH    : integer := 1;
			COMMAND_FIFO_DEPTH  : integer := 4;
			RESPONSE_FIFO_DEPTH : integer := 4;
			MASTER_SYNC_DEPTH   : integer := 2;
			SLAVE_SYNC_DEPTH    : integer := 2
		);
		port (
			m0_clk           : in  std_logic                     := 'X';             -- clk
			m0_reset         : in  std_logic                     := 'X';             -- reset
			s0_clk           : in  std_logic                     := 'X';             -- clk
			s0_reset         : in  std_logic                     := 'X';             -- reset
			s0_waitrequest   : out std_logic;                                        -- waitrequest
			s0_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			s0_readdatavalid : out std_logic;                                        -- readdatavalid
			s0_burstcount    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			s0_address       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			s0_write         : in  std_logic                     := 'X';             -- write
			s0_read          : in  std_logic                     := 'X';             -- read
			s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			s0_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			m0_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			m0_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			m0_burstcount    : out std_logic_vector(0 downto 0);                     -- burstcount
			m0_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			m0_address       : out std_logic_vector(9 downto 0);                     -- address
			m0_write         : out std_logic;                                        -- write
			m0_read          : out std_logic;                                        -- read
			m0_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess   : out std_logic                                         -- debugaccess
		);
	end component altera_avalon_mm_clock_crossing_bridge;

	component nios2_c_tightly_coupled_data_memory is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X'              -- reset_req
		);
	end component nios2_c_tightly_coupled_data_memory;

	component nios2_c_key is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component nios2_c_key;

	component nios2_c_timer_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component nios2_c_timer_0;

	component nios2_c_ledg is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component nios2_c_ledg;

	component nios2_c_to_hex is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(13 downto 0)                     -- export
		);
	end component nios2_c_to_hex;

	component nios2_c_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                                         : in  std_logic                     := 'X';             -- clk
			pll_100_outclk0_clk                                                   : in  std_logic                     := 'X';             -- clk
			cpu_reset_n_reset_bridge_in_reset_reset                               : in  std_logic                     := 'X';             -- reset
			jtag_uart_reset_reset_bridge_in_reset_reset                           : in  std_logic                     := 'X';             -- reset
			mm_clock_crossing_bridge_0_s0_reset_reset_bridge_in_reset_reset       : in  std_logic                     := 'X';             -- reset
			tightly_coupled_instruction_memory_reset2_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			cpu_data_master_address                                               : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			cpu_data_master_waitrequest                                           : out std_logic;                                        -- waitrequest
			cpu_data_master_burstcount                                            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- burstcount
			cpu_data_master_byteenable                                            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_data_master_read                                                  : in  std_logic                     := 'X';             -- read
			cpu_data_master_readdata                                              : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_data_master_readdatavalid                                         : out std_logic;                                        -- readdatavalid
			cpu_data_master_write                                                 : in  std_logic                     := 'X';             -- write
			cpu_data_master_writedata                                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_data_master_debugaccess                                           : in  std_logic                     := 'X';             -- debugaccess
			cpu_instruction_master_address                                        : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address
			cpu_instruction_master_waitrequest                                    : out std_logic;                                        -- waitrequest
			cpu_instruction_master_burstcount                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- burstcount
			cpu_instruction_master_read                                           : in  std_logic                     := 'X';             -- read
			cpu_instruction_master_readdata                                       : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_instruction_master_readdatavalid                                  : out std_logic;                                        -- readdatavalid
			cpu_jtag_debug_module_address                                         : out std_logic_vector(8 downto 0);                     -- address
			cpu_jtag_debug_module_write                                           : out std_logic;                                        -- write
			cpu_jtag_debug_module_read                                            : out std_logic;                                        -- read
			cpu_jtag_debug_module_readdata                                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_jtag_debug_module_writedata                                       : out std_logic_vector(31 downto 0);                    -- writedata
			cpu_jtag_debug_module_byteenable                                      : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_jtag_debug_module_waitrequest                                     : in  std_logic                     := 'X';             -- waitrequest
			cpu_jtag_debug_module_debugaccess                                     : out std_logic;                                        -- debugaccess
			jtag_uart_avalon_jtag_slave_address                                   : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write                                     : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read                                      : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata                                 : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest                               : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                                : out std_logic;                                        -- chipselect
			mm_clock_crossing_bridge_0_s0_address                                 : out std_logic_vector(9 downto 0);                     -- address
			mm_clock_crossing_bridge_0_s0_write                                   : out std_logic;                                        -- write
			mm_clock_crossing_bridge_0_s0_read                                    : out std_logic;                                        -- read
			mm_clock_crossing_bridge_0_s0_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			mm_clock_crossing_bridge_0_s0_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			mm_clock_crossing_bridge_0_s0_burstcount                              : out std_logic_vector(0 downto 0);                     -- burstcount
			mm_clock_crossing_bridge_0_s0_byteenable                              : out std_logic_vector(3 downto 0);                     -- byteenable
			mm_clock_crossing_bridge_0_s0_readdatavalid                           : in  std_logic                     := 'X';             -- readdatavalid
			mm_clock_crossing_bridge_0_s0_waitrequest                             : in  std_logic                     := 'X';             -- waitrequest
			mm_clock_crossing_bridge_0_s0_debugaccess                             : out std_logic;                                        -- debugaccess
			sysid_qsys_0_control_slave_address                                    : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_0_control_slave_readdata                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			tightly_coupled_instruction_memory_s2_address                         : out std_logic_vector(14 downto 0);                    -- address
			tightly_coupled_instruction_memory_s2_write                           : out std_logic;                                        -- write
			tightly_coupled_instruction_memory_s2_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			tightly_coupled_instruction_memory_s2_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			tightly_coupled_instruction_memory_s2_byteenable                      : out std_logic_vector(3 downto 0);                     -- byteenable
			tightly_coupled_instruction_memory_s2_chipselect                      : out std_logic;                                        -- chipselect
			tightly_coupled_instruction_memory_s2_clken                           : out std_logic                                         -- clken
		);
	end component nios2_c_mm_interconnect_0;

	component nios2_c_mm_interconnect_1 is
		port (
			clk_0_clk_clk                                                   : in  std_logic                     := 'X';             -- clk
			key_reset_reset_bridge_in_reset_reset                           : in  std_logic                     := 'X';             -- reset
			mm_clock_crossing_bridge_0_m0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			mm_clock_crossing_bridge_0_m0_address                           : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			mm_clock_crossing_bridge_0_m0_waitrequest                       : out std_logic;                                        -- waitrequest
			mm_clock_crossing_bridge_0_m0_burstcount                        : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			mm_clock_crossing_bridge_0_m0_byteenable                        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			mm_clock_crossing_bridge_0_m0_read                              : in  std_logic                     := 'X';             -- read
			mm_clock_crossing_bridge_0_m0_readdata                          : out std_logic_vector(31 downto 0);                    -- readdata
			mm_clock_crossing_bridge_0_m0_readdatavalid                     : out std_logic;                                        -- readdatavalid
			mm_clock_crossing_bridge_0_m0_write                             : in  std_logic                     := 'X';             -- write
			mm_clock_crossing_bridge_0_m0_writedata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			mm_clock_crossing_bridge_0_m0_debugaccess                       : in  std_logic                     := 'X';             -- debugaccess
			key_s1_address                                                  : out std_logic_vector(1 downto 0);                     -- address
			key_s1_write                                                    : out std_logic;                                        -- write
			key_s1_readdata                                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			key_s1_writedata                                                : out std_logic_vector(31 downto 0);                    -- writedata
			key_s1_chipselect                                               : out std_logic;                                        -- chipselect
			ledg_s1_address                                                 : out std_logic_vector(1 downto 0);                     -- address
			ledg_s1_write                                                   : out std_logic;                                        -- write
			ledg_s1_readdata                                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			ledg_s1_writedata                                               : out std_logic_vector(31 downto 0);                    -- writedata
			ledg_s1_chipselect                                              : out std_logic;                                        -- chipselect
			timer_0_s1_address                                              : out std_logic_vector(2 downto 0);                     -- address
			timer_0_s1_write                                                : out std_logic;                                        -- write
			timer_0_s1_readdata                                             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_0_s1_writedata                                            : out std_logic_vector(15 downto 0);                    -- writedata
			timer_0_s1_chipselect                                           : out std_logic;                                        -- chipselect
			to_hex_s1_address                                               : out std_logic_vector(1 downto 0);                     -- address
			to_hex_s1_write                                                 : out std_logic;                                        -- write
			to_hex_s1_readdata                                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			to_hex_s1_writedata                                             : out std_logic_vector(31 downto 0);                    -- writedata
			to_hex_s1_chipselect                                            : out std_logic                                         -- chipselect
		);
	end component nios2_c_mm_interconnect_1;

	component nios2_c_mm_interconnect_2 is
		port (
			clk_0_clk_clk                                          : in  std_logic                     := 'X';             -- clk
			cpu_reset_n_reset_bridge_in_reset_reset                : in  std_logic                     := 'X';             -- reset
			cpu_tightly_coupled_instruction_master_0_address       : in  std_logic_vector(16 downto 0) := (others => 'X'); -- address
			cpu_tightly_coupled_instruction_master_0_waitrequest   : out std_logic;                                        -- waitrequest
			cpu_tightly_coupled_instruction_master_0_read          : in  std_logic                     := 'X';             -- read
			cpu_tightly_coupled_instruction_master_0_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_tightly_coupled_instruction_master_0_readdatavalid : out std_logic;                                        -- readdatavalid
			cpu_tightly_coupled_instruction_master_0_clken         : in  std_logic                     := 'X';             -- clken
			tightly_coupled_instruction_memory_s1_address          : out std_logic_vector(14 downto 0);                    -- address
			tightly_coupled_instruction_memory_s1_write            : out std_logic;                                        -- write
			tightly_coupled_instruction_memory_s1_readdata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			tightly_coupled_instruction_memory_s1_writedata        : out std_logic_vector(31 downto 0);                    -- writedata
			tightly_coupled_instruction_memory_s1_byteenable       : out std_logic_vector(3 downto 0);                     -- byteenable
			tightly_coupled_instruction_memory_s1_chipselect       : out std_logic;                                        -- chipselect
			tightly_coupled_instruction_memory_s1_clken            : out std_logic                                         -- clken
		);
	end component nios2_c_mm_interconnect_2;

	component nios2_c_mm_interconnect_3 is
		port (
			clk_0_clk_clk                                   : in  std_logic                     := 'X';             -- clk
			cpu_reset_n_reset_bridge_in_reset_reset         : in  std_logic                     := 'X';             -- reset
			cpu_tightly_coupled_data_master_0_address       : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address
			cpu_tightly_coupled_data_master_0_waitrequest   : out std_logic;                                        -- waitrequest
			cpu_tightly_coupled_data_master_0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_tightly_coupled_data_master_0_read          : in  std_logic                     := 'X';             -- read
			cpu_tightly_coupled_data_master_0_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_tightly_coupled_data_master_0_readdatavalid : out std_logic;                                        -- readdatavalid
			cpu_tightly_coupled_data_master_0_write         : in  std_logic                     := 'X';             -- write
			cpu_tightly_coupled_data_master_0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_tightly_coupled_data_master_0_clken         : in  std_logic                     := 'X';             -- clken
			tightly_coupled_data_memory_s1_address          : out std_logic_vector(12 downto 0);                    -- address
			tightly_coupled_data_memory_s1_write            : out std_logic;                                        -- write
			tightly_coupled_data_memory_s1_readdata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			tightly_coupled_data_memory_s1_writedata        : out std_logic_vector(31 downto 0);                    -- writedata
			tightly_coupled_data_memory_s1_byteenable       : out std_logic_vector(3 downto 0);                     -- byteenable
			tightly_coupled_data_memory_s1_chipselect       : out std_logic;                                        -- chipselect
			tightly_coupled_data_memory_s1_clken            : out std_logic                                         -- clken
		);
	end component nios2_c_mm_interconnect_3;

	component nios2_c_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component nios2_c_irq_mapper;

	component altera_irq_clock_crosser is
		generic (
			IRQ_WIDTH : integer := 1
		);
		port (
			receiver_clk   : in  std_logic                    := 'X';             -- clk
			sender_clk     : in  std_logic                    := 'X';             -- clk
			receiver_reset : in  std_logic                    := 'X';             -- reset
			sender_reset   : in  std_logic                    := 'X';             -- reset
			receiver_irq   : in  std_logic_vector(0 downto 0) := (others => 'X'); -- irq
			sender_irq     : out std_logic_vector(0 downto 0)                     -- irq
		);
	end component altera_irq_clock_crosser;

	component nios2_c_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component nios2_c_rst_controller;

	component nios2_c_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component nios2_c_rst_controller_001;

	component nios2_c_rst_controller_002 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component nios2_c_rst_controller_002;

	component nios2_c_rst_controller_003 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component nios2_c_rst_controller_003;

	signal pll_100_outclk0_clk                                                : std_logic;                     -- pll_100:outclk_0 -> [irq_synchronizer:receiver_clk, jtag_uart:clk, mm_clock_crossing_bridge_0:s0_clk, mm_interconnect_0:pll_100_outclk0_clk, rst_controller_002:clk, rst_controller_003:clk]
	signal mm_interconnect_0_mm_clock_crossing_bridge_0_s0_waitrequest        : std_logic;                     -- mm_clock_crossing_bridge_0:s0_waitrequest -> mm_interconnect_0:mm_clock_crossing_bridge_0_s0_waitrequest
	signal mm_interconnect_0_mm_clock_crossing_bridge_0_s0_burstcount         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:mm_clock_crossing_bridge_0_s0_burstcount -> mm_clock_crossing_bridge_0:s0_burstcount
	signal mm_interconnect_0_mm_clock_crossing_bridge_0_s0_writedata          : std_logic_vector(31 downto 0); -- mm_interconnect_0:mm_clock_crossing_bridge_0_s0_writedata -> mm_clock_crossing_bridge_0:s0_writedata
	signal mm_interconnect_0_mm_clock_crossing_bridge_0_s0_address            : std_logic_vector(9 downto 0);  -- mm_interconnect_0:mm_clock_crossing_bridge_0_s0_address -> mm_clock_crossing_bridge_0:s0_address
	signal mm_interconnect_0_mm_clock_crossing_bridge_0_s0_write              : std_logic;                     -- mm_interconnect_0:mm_clock_crossing_bridge_0_s0_write -> mm_clock_crossing_bridge_0:s0_write
	signal mm_interconnect_0_mm_clock_crossing_bridge_0_s0_read               : std_logic;                     -- mm_interconnect_0:mm_clock_crossing_bridge_0_s0_read -> mm_clock_crossing_bridge_0:s0_read
	signal mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdata           : std_logic_vector(31 downto 0); -- mm_clock_crossing_bridge_0:s0_readdata -> mm_interconnect_0:mm_clock_crossing_bridge_0_s0_readdata
	signal mm_interconnect_0_mm_clock_crossing_bridge_0_s0_debugaccess        : std_logic;                     -- mm_interconnect_0:mm_clock_crossing_bridge_0_s0_debugaccess -> mm_clock_crossing_bridge_0:s0_debugaccess
	signal mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdatavalid      : std_logic;                     -- mm_clock_crossing_bridge_0:s0_readdatavalid -> mm_interconnect_0:mm_clock_crossing_bridge_0_s0_readdatavalid
	signal mm_interconnect_0_mm_clock_crossing_bridge_0_s0_byteenable         : std_logic_vector(3 downto 0);  -- mm_interconnect_0:mm_clock_crossing_bridge_0_s0_byteenable -> mm_clock_crossing_bridge_0:s0_byteenable
	signal cpu_instruction_master_burstcount                                  : std_logic_vector(3 downto 0);  -- cpu:i_burstcount -> mm_interconnect_0:cpu_instruction_master_burstcount
	signal cpu_instruction_master_waitrequest                                 : std_logic;                     -- mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	signal cpu_instruction_master_address                                     : std_logic_vector(18 downto 0); -- cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	signal cpu_instruction_master_read                                        : std_logic;                     -- cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	signal cpu_instruction_master_readdata                                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	signal cpu_instruction_master_readdatavalid                               : std_logic;                     -- mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	signal mm_interconnect_0_cpu_jtag_debug_module_waitrequest                : std_logic;                     -- cpu:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_jtag_debug_module_waitrequest
	signal mm_interconnect_0_cpu_jtag_debug_module_writedata                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_jtag_debug_module_writedata -> cpu:jtag_debug_module_writedata
	signal mm_interconnect_0_cpu_jtag_debug_module_address                    : std_logic_vector(8 downto 0);  -- mm_interconnect_0:cpu_jtag_debug_module_address -> cpu:jtag_debug_module_address
	signal mm_interconnect_0_cpu_jtag_debug_module_write                      : std_logic;                     -- mm_interconnect_0:cpu_jtag_debug_module_write -> cpu:jtag_debug_module_write
	signal mm_interconnect_0_cpu_jtag_debug_module_read                       : std_logic;                     -- mm_interconnect_0:cpu_jtag_debug_module_read -> cpu:jtag_debug_module_read
	signal mm_interconnect_0_cpu_jtag_debug_module_readdata                   : std_logic_vector(31 downto 0); -- cpu:jtag_debug_module_readdata -> mm_interconnect_0:cpu_jtag_debug_module_readdata
	signal mm_interconnect_0_cpu_jtag_debug_module_debugaccess                : std_logic;                     -- mm_interconnect_0:cpu_jtag_debug_module_debugaccess -> cpu:jtag_debug_module_debugaccess
	signal mm_interconnect_0_cpu_jtag_debug_module_byteenable                 : std_logic_vector(3 downto 0);  -- mm_interconnect_0:cpu_jtag_debug_module_byteenable -> cpu:jtag_debug_module_byteenable
	signal mm_interconnect_0_tightly_coupled_instruction_memory_s2_writedata  : std_logic_vector(31 downto 0); -- mm_interconnect_0:tightly_coupled_instruction_memory_s2_writedata -> tightly_coupled_instruction_memory:writedata2
	signal mm_interconnect_0_tightly_coupled_instruction_memory_s2_address    : std_logic_vector(14 downto 0); -- mm_interconnect_0:tightly_coupled_instruction_memory_s2_address -> tightly_coupled_instruction_memory:address2
	signal mm_interconnect_0_tightly_coupled_instruction_memory_s2_chipselect : std_logic;                     -- mm_interconnect_0:tightly_coupled_instruction_memory_s2_chipselect -> tightly_coupled_instruction_memory:chipselect2
	signal mm_interconnect_0_tightly_coupled_instruction_memory_s2_clken      : std_logic;                     -- mm_interconnect_0:tightly_coupled_instruction_memory_s2_clken -> tightly_coupled_instruction_memory:clken2
	signal mm_interconnect_0_tightly_coupled_instruction_memory_s2_write      : std_logic;                     -- mm_interconnect_0:tightly_coupled_instruction_memory_s2_write -> tightly_coupled_instruction_memory:write2
	signal mm_interconnect_0_tightly_coupled_instruction_memory_s2_readdata   : std_logic_vector(31 downto 0); -- tightly_coupled_instruction_memory:readdata2 -> mm_interconnect_0:tightly_coupled_instruction_memory_s2_readdata
	signal mm_interconnect_0_tightly_coupled_instruction_memory_s2_byteenable : std_logic_vector(3 downto 0);  -- mm_interconnect_0:tightly_coupled_instruction_memory_s2_byteenable -> tightly_coupled_instruction_memory:byteenable2
	signal mm_interconnect_0_sysid_qsys_0_control_slave_address               : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	signal mm_interconnect_0_sysid_qsys_0_control_slave_readdata              : std_logic_vector(31 downto 0); -- sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest          : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata            : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address              : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect           : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write                : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read                 : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata             : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	signal cpu_data_master_burstcount                                         : std_logic_vector(3 downto 0);  -- cpu:d_burstcount -> mm_interconnect_0:cpu_data_master_burstcount
	signal cpu_data_master_waitrequest                                        : std_logic;                     -- mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	signal cpu_data_master_writedata                                          : std_logic_vector(31 downto 0); -- cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	signal cpu_data_master_address                                            : std_logic_vector(24 downto 0); -- cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	signal cpu_data_master_write                                              : std_logic;                     -- cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	signal cpu_data_master_read                                               : std_logic;                     -- cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	signal cpu_data_master_readdata                                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	signal cpu_data_master_debugaccess                                        : std_logic;                     -- cpu:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	signal cpu_data_master_readdatavalid                                      : std_logic;                     -- mm_interconnect_0:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	signal cpu_data_master_byteenable                                         : std_logic_vector(3 downto 0);  -- cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	signal mm_interconnect_1_to_hex_s1_writedata                              : std_logic_vector(31 downto 0); -- mm_interconnect_1:to_hex_s1_writedata -> to_hex:writedata
	signal mm_interconnect_1_to_hex_s1_address                                : std_logic_vector(1 downto 0);  -- mm_interconnect_1:to_hex_s1_address -> to_hex:address
	signal mm_interconnect_1_to_hex_s1_chipselect                             : std_logic;                     -- mm_interconnect_1:to_hex_s1_chipselect -> to_hex:chipselect
	signal mm_interconnect_1_to_hex_s1_write                                  : std_logic;                     -- mm_interconnect_1:to_hex_s1_write -> mm_interconnect_1_to_hex_s1_write:in
	signal mm_interconnect_1_to_hex_s1_readdata                               : std_logic_vector(31 downto 0); -- to_hex:readdata -> mm_interconnect_1:to_hex_s1_readdata
	signal mm_interconnect_1_key_s1_writedata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_1:key_s1_writedata -> key:writedata
	signal mm_interconnect_1_key_s1_address                                   : std_logic_vector(1 downto 0);  -- mm_interconnect_1:key_s1_address -> key:address
	signal mm_interconnect_1_key_s1_chipselect                                : std_logic;                     -- mm_interconnect_1:key_s1_chipselect -> key:chipselect
	signal mm_interconnect_1_key_s1_write                                     : std_logic;                     -- mm_interconnect_1:key_s1_write -> mm_interconnect_1_key_s1_write:in
	signal mm_interconnect_1_key_s1_readdata                                  : std_logic_vector(31 downto 0); -- key:readdata -> mm_interconnect_1:key_s1_readdata
	signal mm_clock_crossing_bridge_0_m0_burstcount                           : std_logic_vector(0 downto 0);  -- mm_clock_crossing_bridge_0:m0_burstcount -> mm_interconnect_1:mm_clock_crossing_bridge_0_m0_burstcount
	signal mm_clock_crossing_bridge_0_m0_waitrequest                          : std_logic;                     -- mm_interconnect_1:mm_clock_crossing_bridge_0_m0_waitrequest -> mm_clock_crossing_bridge_0:m0_waitrequest
	signal mm_clock_crossing_bridge_0_m0_address                              : std_logic_vector(9 downto 0);  -- mm_clock_crossing_bridge_0:m0_address -> mm_interconnect_1:mm_clock_crossing_bridge_0_m0_address
	signal mm_clock_crossing_bridge_0_m0_writedata                            : std_logic_vector(31 downto 0); -- mm_clock_crossing_bridge_0:m0_writedata -> mm_interconnect_1:mm_clock_crossing_bridge_0_m0_writedata
	signal mm_clock_crossing_bridge_0_m0_write                                : std_logic;                     -- mm_clock_crossing_bridge_0:m0_write -> mm_interconnect_1:mm_clock_crossing_bridge_0_m0_write
	signal mm_clock_crossing_bridge_0_m0_read                                 : std_logic;                     -- mm_clock_crossing_bridge_0:m0_read -> mm_interconnect_1:mm_clock_crossing_bridge_0_m0_read
	signal mm_clock_crossing_bridge_0_m0_readdata                             : std_logic_vector(31 downto 0); -- mm_interconnect_1:mm_clock_crossing_bridge_0_m0_readdata -> mm_clock_crossing_bridge_0:m0_readdata
	signal mm_clock_crossing_bridge_0_m0_debugaccess                          : std_logic;                     -- mm_clock_crossing_bridge_0:m0_debugaccess -> mm_interconnect_1:mm_clock_crossing_bridge_0_m0_debugaccess
	signal mm_clock_crossing_bridge_0_m0_byteenable                           : std_logic_vector(3 downto 0);  -- mm_clock_crossing_bridge_0:m0_byteenable -> mm_interconnect_1:mm_clock_crossing_bridge_0_m0_byteenable
	signal mm_clock_crossing_bridge_0_m0_readdatavalid                        : std_logic;                     -- mm_interconnect_1:mm_clock_crossing_bridge_0_m0_readdatavalid -> mm_clock_crossing_bridge_0:m0_readdatavalid
	signal mm_interconnect_1_ledg_s1_writedata                                : std_logic_vector(31 downto 0); -- mm_interconnect_1:ledg_s1_writedata -> ledg:writedata
	signal mm_interconnect_1_ledg_s1_address                                  : std_logic_vector(1 downto 0);  -- mm_interconnect_1:ledg_s1_address -> ledg:address
	signal mm_interconnect_1_ledg_s1_chipselect                               : std_logic;                     -- mm_interconnect_1:ledg_s1_chipselect -> ledg:chipselect
	signal mm_interconnect_1_ledg_s1_write                                    : std_logic;                     -- mm_interconnect_1:ledg_s1_write -> mm_interconnect_1_ledg_s1_write:in
	signal mm_interconnect_1_ledg_s1_readdata                                 : std_logic_vector(31 downto 0); -- ledg:readdata -> mm_interconnect_1:ledg_s1_readdata
	signal mm_interconnect_1_timer_0_s1_writedata                             : std_logic_vector(15 downto 0); -- mm_interconnect_1:timer_0_s1_writedata -> timer_0:writedata
	signal mm_interconnect_1_timer_0_s1_address                               : std_logic_vector(2 downto 0);  -- mm_interconnect_1:timer_0_s1_address -> timer_0:address
	signal mm_interconnect_1_timer_0_s1_chipselect                            : std_logic;                     -- mm_interconnect_1:timer_0_s1_chipselect -> timer_0:chipselect
	signal mm_interconnect_1_timer_0_s1_write                                 : std_logic;                     -- mm_interconnect_1:timer_0_s1_write -> mm_interconnect_1_timer_0_s1_write:in
	signal mm_interconnect_1_timer_0_s1_readdata                              : std_logic_vector(15 downto 0); -- timer_0:readdata -> mm_interconnect_1:timer_0_s1_readdata
	signal mm_interconnect_2_tightly_coupled_instruction_memory_s1_writedata  : std_logic_vector(31 downto 0); -- mm_interconnect_2:tightly_coupled_instruction_memory_s1_writedata -> tightly_coupled_instruction_memory:writedata
	signal mm_interconnect_2_tightly_coupled_instruction_memory_s1_address    : std_logic_vector(14 downto 0); -- mm_interconnect_2:tightly_coupled_instruction_memory_s1_address -> tightly_coupled_instruction_memory:address
	signal mm_interconnect_2_tightly_coupled_instruction_memory_s1_chipselect : std_logic;                     -- mm_interconnect_2:tightly_coupled_instruction_memory_s1_chipselect -> tightly_coupled_instruction_memory:chipselect
	signal mm_interconnect_2_tightly_coupled_instruction_memory_s1_clken      : std_logic;                     -- mm_interconnect_2:tightly_coupled_instruction_memory_s1_clken -> tightly_coupled_instruction_memory:clken
	signal mm_interconnect_2_tightly_coupled_instruction_memory_s1_write      : std_logic;                     -- mm_interconnect_2:tightly_coupled_instruction_memory_s1_write -> tightly_coupled_instruction_memory:write
	signal mm_interconnect_2_tightly_coupled_instruction_memory_s1_readdata   : std_logic_vector(31 downto 0); -- tightly_coupled_instruction_memory:readdata -> mm_interconnect_2:tightly_coupled_instruction_memory_s1_readdata
	signal mm_interconnect_2_tightly_coupled_instruction_memory_s1_byteenable : std_logic_vector(3 downto 0);  -- mm_interconnect_2:tightly_coupled_instruction_memory_s1_byteenable -> tightly_coupled_instruction_memory:byteenable
	signal cpu_tightly_coupled_instruction_master_0_waitrequest               : std_logic;                     -- mm_interconnect_2:cpu_tightly_coupled_instruction_master_0_waitrequest -> cpu:icm0_waitrequest
	signal cpu_tightly_coupled_instruction_master_0_address                   : std_logic_vector(16 downto 0); -- cpu:icm0_address -> mm_interconnect_2:cpu_tightly_coupled_instruction_master_0_address
	signal cpu_tightly_coupled_instruction_master_0_clken                     : std_logic;                     -- cpu:icm0_clken -> mm_interconnect_2:cpu_tightly_coupled_instruction_master_0_clken
	signal cpu_tightly_coupled_instruction_master_0_read                      : std_logic;                     -- cpu:icm0_read -> mm_interconnect_2:cpu_tightly_coupled_instruction_master_0_read
	signal cpu_tightly_coupled_instruction_master_0_readdata                  : std_logic_vector(31 downto 0); -- mm_interconnect_2:cpu_tightly_coupled_instruction_master_0_readdata -> cpu:icm0_readdata
	signal cpu_tightly_coupled_instruction_master_0_readdatavalid             : std_logic;                     -- mm_interconnect_2:cpu_tightly_coupled_instruction_master_0_readdatavalid -> cpu:icm0_readdatavalid
	signal mm_interconnect_3_tightly_coupled_data_memory_s1_writedata         : std_logic_vector(31 downto 0); -- mm_interconnect_3:tightly_coupled_data_memory_s1_writedata -> tightly_coupled_data_memory:writedata
	signal mm_interconnect_3_tightly_coupled_data_memory_s1_address           : std_logic_vector(12 downto 0); -- mm_interconnect_3:tightly_coupled_data_memory_s1_address -> tightly_coupled_data_memory:address
	signal mm_interconnect_3_tightly_coupled_data_memory_s1_chipselect        : std_logic;                     -- mm_interconnect_3:tightly_coupled_data_memory_s1_chipselect -> tightly_coupled_data_memory:chipselect
	signal mm_interconnect_3_tightly_coupled_data_memory_s1_clken             : std_logic;                     -- mm_interconnect_3:tightly_coupled_data_memory_s1_clken -> tightly_coupled_data_memory:clken
	signal mm_interconnect_3_tightly_coupled_data_memory_s1_write             : std_logic;                     -- mm_interconnect_3:tightly_coupled_data_memory_s1_write -> tightly_coupled_data_memory:write
	signal mm_interconnect_3_tightly_coupled_data_memory_s1_readdata          : std_logic_vector(31 downto 0); -- tightly_coupled_data_memory:readdata -> mm_interconnect_3:tightly_coupled_data_memory_s1_readdata
	signal mm_interconnect_3_tightly_coupled_data_memory_s1_byteenable        : std_logic_vector(3 downto 0);  -- mm_interconnect_3:tightly_coupled_data_memory_s1_byteenable -> tightly_coupled_data_memory:byteenable
	signal cpu_tightly_coupled_data_master_0_waitrequest                      : std_logic;                     -- mm_interconnect_3:cpu_tightly_coupled_data_master_0_waitrequest -> cpu:dcm0_waitrequest
	signal cpu_tightly_coupled_data_master_0_writedata                        : std_logic_vector(31 downto 0); -- cpu:dcm0_writedata -> mm_interconnect_3:cpu_tightly_coupled_data_master_0_writedata
	signal cpu_tightly_coupled_data_master_0_address                          : std_logic_vector(18 downto 0); -- cpu:dcm0_address -> mm_interconnect_3:cpu_tightly_coupled_data_master_0_address
	signal cpu_tightly_coupled_data_master_0_clken                            : std_logic;                     -- cpu:dcm0_clken -> mm_interconnect_3:cpu_tightly_coupled_data_master_0_clken
	signal cpu_tightly_coupled_data_master_0_write                            : std_logic;                     -- cpu:dcm0_write -> mm_interconnect_3:cpu_tightly_coupled_data_master_0_write
	signal cpu_tightly_coupled_data_master_0_read                             : std_logic;                     -- cpu:dcm0_read -> mm_interconnect_3:cpu_tightly_coupled_data_master_0_read
	signal cpu_tightly_coupled_data_master_0_readdata                         : std_logic_vector(31 downto 0); -- mm_interconnect_3:cpu_tightly_coupled_data_master_0_readdata -> cpu:dcm0_readdata
	signal cpu_tightly_coupled_data_master_0_byteenable                       : std_logic_vector(3 downto 0);  -- cpu:dcm0_byteenable -> mm_interconnect_3:cpu_tightly_coupled_data_master_0_byteenable
	signal cpu_tightly_coupled_data_master_0_readdatavalid                    : std_logic;                     -- mm_interconnect_3:cpu_tightly_coupled_data_master_0_readdatavalid -> cpu:dcm0_readdatavalid
	signal irq_mapper_receiver1_irq                                           : std_logic;                     -- key:irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                           : std_logic;                     -- timer_0:irq -> irq_mapper:receiver2_irq
	signal cpu_d_irq_irq                                                      : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> cpu:d_irq
	signal irq_mapper_receiver0_irq                                           : std_logic;                     -- irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	signal irq_synchronizer_receiver_irq                                      : std_logic_vector(0 downto 0);  -- jtag_uart:av_irq -> irq_synchronizer:receiver_irq
	signal rst_controller_reset_out_reset                                     : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, irq_synchronizer:sender_reset, mm_clock_crossing_bridge_0:m0_reset, mm_interconnect_0:cpu_reset_n_reset_bridge_in_reset_reset, mm_interconnect_1:mm_clock_crossing_bridge_0_m0_reset_reset_bridge_in_reset_reset, mm_interconnect_2:cpu_reset_n_reset_bridge_in_reset_reset, mm_interconnect_3:cpu_reset_n_reset_bridge_in_reset_reset, pll_100:rst, rst_controller_reset_out_reset:in, rst_translator:in_reset, tightly_coupled_data_memory:reset, tightly_coupled_instruction_memory:reset]
	signal rst_controller_reset_out_reset_req                                 : std_logic;                     -- rst_controller:reset_req -> [cpu:reset_req, rst_translator:reset_req_in, tightly_coupled_data_memory:reset_req, tightly_coupled_instruction_memory:reset_req]
	signal cpu_jtag_debug_module_reset_reset                                  : std_logic;                     -- cpu:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_002:reset_in1]
	signal rst_controller_001_reset_out_reset                                 : std_logic;                     -- rst_controller_001:reset_out -> [mm_interconnect_0:tightly_coupled_instruction_memory_reset2_reset_bridge_in_reset_reset, mm_interconnect_1:key_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in, rst_translator_001:in_reset, tightly_coupled_instruction_memory:reset2]
	signal rst_controller_001_reset_out_reset_req                             : std_logic;                     -- rst_controller_001:reset_req -> [rst_translator_001:reset_req_in, tightly_coupled_instruction_memory:reset_req2]
	signal rst_controller_002_reset_out_reset                                 : std_logic;                     -- rst_controller_002:reset_out -> [irq_synchronizer:receiver_reset, mm_interconnect_0:jtag_uart_reset_reset_bridge_in_reset_reset, rst_controller_002_reset_out_reset:in]
	signal rst_controller_003_reset_out_reset                                 : std_logic;                     -- rst_controller_003:reset_out -> [mm_clock_crossing_bridge_0:s0_reset, mm_interconnect_0:mm_clock_crossing_bridge_0_s0_reset_reset_bridge_in_reset_reset]
	signal reset_reset_n_ports_inv                                            : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0, rst_controller_003:reset_in0]
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv      : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv       : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_1_to_hex_s1_write_ports_inv                        : std_logic;                     -- mm_interconnect_1_to_hex_s1_write:inv -> to_hex:write_n
	signal mm_interconnect_1_key_s1_write_ports_inv                           : std_logic;                     -- mm_interconnect_1_key_s1_write:inv -> key:write_n
	signal mm_interconnect_1_ledg_s1_write_ports_inv                          : std_logic;                     -- mm_interconnect_1_ledg_s1_write:inv -> ledg:write_n
	signal mm_interconnect_1_timer_0_s1_write_ports_inv                       : std_logic;                     -- mm_interconnect_1_timer_0_s1_write:inv -> timer_0:write_n
	signal rst_controller_reset_out_reset_ports_inv                           : std_logic;                     -- rst_controller_reset_out_reset:inv -> [cpu:reset_n, sysid_qsys_0:reset_n]
	signal rst_controller_001_reset_out_reset_ports_inv                       : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> [key:reset_n, ledg:reset_n, timer_0:reset_n, to_hex:reset_n]
	signal rst_controller_002_reset_out_reset_ports_inv                       : std_logic;                     -- rst_controller_002_reset_out_reset:inv -> jtag_uart:rst_n

begin

	cpu : component nios2_c_cpu
		port map (
			clk                                   => clk_clk,                                                --                                  clk.clk
			reset_n                               => rst_controller_reset_out_reset_ports_inv,               --                              reset_n.reset_n
			reset_req                             => rst_controller_reset_out_reset_req,                     --                                     .reset_req
			d_address                             => cpu_data_master_address,                                --                          data_master.address
			d_byteenable                          => cpu_data_master_byteenable,                             --                                     .byteenable
			d_read                                => cpu_data_master_read,                                   --                                     .read
			d_readdata                            => cpu_data_master_readdata,                               --                                     .readdata
			d_waitrequest                         => cpu_data_master_waitrequest,                            --                                     .waitrequest
			d_write                               => cpu_data_master_write,                                  --                                     .write
			d_writedata                           => cpu_data_master_writedata,                              --                                     .writedata
			d_burstcount                          => cpu_data_master_burstcount,                             --                                     .burstcount
			d_readdatavalid                       => cpu_data_master_readdatavalid,                          --                                     .readdatavalid
			jtag_debug_module_debugaccess_to_roms => cpu_data_master_debugaccess,                            --                                     .debugaccess
			i_address                             => cpu_instruction_master_address,                         --                   instruction_master.address
			i_read                                => cpu_instruction_master_read,                            --                                     .read
			i_readdata                            => cpu_instruction_master_readdata,                        --                                     .readdata
			i_waitrequest                         => cpu_instruction_master_waitrequest,                     --                                     .waitrequest
			i_burstcount                          => cpu_instruction_master_burstcount,                      --                                     .burstcount
			i_readdatavalid                       => cpu_instruction_master_readdatavalid,                   --                                     .readdatavalid
			dcm0_readdata                         => cpu_tightly_coupled_data_master_0_readdata,             --        tightly_coupled_data_master_0.readdata
			dcm0_waitrequest                      => cpu_tightly_coupled_data_master_0_waitrequest,          --                                     .waitrequest
			dcm0_readdatavalid                    => cpu_tightly_coupled_data_master_0_readdatavalid,        --                                     .readdatavalid
			dcm0_address                          => cpu_tightly_coupled_data_master_0_address,              --                                     .address
			dcm0_read                             => cpu_tightly_coupled_data_master_0_read,                 --                                     .read
			dcm0_clken                            => cpu_tightly_coupled_data_master_0_clken,                --                                     .clken
			dcm0_write                            => cpu_tightly_coupled_data_master_0_write,                --                                     .write
			dcm0_writedata                        => cpu_tightly_coupled_data_master_0_writedata,            --                                     .writedata
			dcm0_byteenable                       => cpu_tightly_coupled_data_master_0_byteenable,           --                                     .byteenable
			icm0_readdata                         => cpu_tightly_coupled_instruction_master_0_readdata,      -- tightly_coupled_instruction_master_0.readdata
			icm0_waitrequest                      => cpu_tightly_coupled_instruction_master_0_waitrequest,   --                                     .waitrequest
			icm0_readdatavalid                    => cpu_tightly_coupled_instruction_master_0_readdatavalid, --                                     .readdatavalid
			icm0_address                          => cpu_tightly_coupled_instruction_master_0_address,       --                                     .address
			icm0_read                             => cpu_tightly_coupled_instruction_master_0_read,          --                                     .read
			icm0_clken                            => cpu_tightly_coupled_instruction_master_0_clken,         --                                     .clken
			d_irq                                 => cpu_d_irq_irq,                                          --                                d_irq.irq
			jtag_debug_module_resetrequest        => cpu_jtag_debug_module_reset_reset,                      --              jtag_debug_module_reset.reset
			jtag_debug_module_address             => mm_interconnect_0_cpu_jtag_debug_module_address,        --                    jtag_debug_module.address
			jtag_debug_module_byteenable          => mm_interconnect_0_cpu_jtag_debug_module_byteenable,     --                                     .byteenable
			jtag_debug_module_debugaccess         => mm_interconnect_0_cpu_jtag_debug_module_debugaccess,    --                                     .debugaccess
			jtag_debug_module_read                => mm_interconnect_0_cpu_jtag_debug_module_read,           --                                     .read
			jtag_debug_module_readdata            => mm_interconnect_0_cpu_jtag_debug_module_readdata,       --                                     .readdata
			jtag_debug_module_waitrequest         => mm_interconnect_0_cpu_jtag_debug_module_waitrequest,    --                                     .waitrequest
			jtag_debug_module_write               => mm_interconnect_0_cpu_jtag_debug_module_write,          --                                     .write
			jtag_debug_module_writedata           => mm_interconnect_0_cpu_jtag_debug_module_writedata,      --                                     .writedata
			no_ci_readra                          => open                                                    --            custom_instruction_master.readra
		);

	tightly_coupled_instruction_memory : component nios2_c_tightly_coupled_instruction_memory
		port map (
			clk         => clk_clk,                                                            --   clk1.clk
			address     => mm_interconnect_2_tightly_coupled_instruction_memory_s1_address,    --     s1.address
			clken       => mm_interconnect_2_tightly_coupled_instruction_memory_s1_clken,      --       .clken
			chipselect  => mm_interconnect_2_tightly_coupled_instruction_memory_s1_chipselect, --       .chipselect
			write       => mm_interconnect_2_tightly_coupled_instruction_memory_s1_write,      --       .write
			readdata    => mm_interconnect_2_tightly_coupled_instruction_memory_s1_readdata,   --       .readdata
			writedata   => mm_interconnect_2_tightly_coupled_instruction_memory_s1_writedata,  --       .writedata
			byteenable  => mm_interconnect_2_tightly_coupled_instruction_memory_s1_byteenable, --       .byteenable
			reset       => rst_controller_reset_out_reset,                                     -- reset1.reset
			reset_req   => rst_controller_reset_out_reset_req,                                 --       .reset_req
			address2    => mm_interconnect_0_tightly_coupled_instruction_memory_s2_address,    --     s2.address
			chipselect2 => mm_interconnect_0_tightly_coupled_instruction_memory_s2_chipselect, --       .chipselect
			clken2      => mm_interconnect_0_tightly_coupled_instruction_memory_s2_clken,      --       .clken
			write2      => mm_interconnect_0_tightly_coupled_instruction_memory_s2_write,      --       .write
			readdata2   => mm_interconnect_0_tightly_coupled_instruction_memory_s2_readdata,   --       .readdata
			writedata2  => mm_interconnect_0_tightly_coupled_instruction_memory_s2_writedata,  --       .writedata
			byteenable2 => mm_interconnect_0_tightly_coupled_instruction_memory_s2_byteenable, --       .byteenable
			clk2        => clk_clk,                                                            --   clk2.clk
			reset2      => rst_controller_001_reset_out_reset,                                 -- reset2.reset
			reset_req2  => rst_controller_001_reset_out_reset_req                              --       .reset_req
		);

	pll_100 : component nios2_c_pll_100
		port map (
			refclk   => clk_clk,                        --  refclk.clk
			rst      => rst_controller_reset_out_reset, --   reset.reset
			outclk_0 => pll_100_outclk0_clk,            -- outclk0.clk
			locked   => open                            -- (terminated)
		);

	jtag_uart : component nios2_c_jtag_uart
		port map (
			clk            => pll_100_outclk0_clk,                                           --               clk.clk
			rst_n          => rst_controller_002_reset_out_reset_ports_inv,                  --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_synchronizer_receiver_irq(0)                               --               irq.irq
		);

	sysid_qsys_0 : component nios2_c_sysid_qsys_0
		port map (
			clock    => clk_clk,                                                 --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,                --         reset.reset_n
			readdata => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_qsys_0_control_slave_address(0)  --              .address
		);

	mm_clock_crossing_bridge_0 : component altera_avalon_mm_clock_crossing_bridge
		generic map (
			DATA_WIDTH          => 32,
			SYMBOL_WIDTH        => 8,
			ADDRESS_WIDTH       => 10,
			BURSTCOUNT_WIDTH    => 1,
			COMMAND_FIFO_DEPTH  => 4,
			RESPONSE_FIFO_DEPTH => 4,
			MASTER_SYNC_DEPTH   => 2,
			SLAVE_SYNC_DEPTH    => 2
		)
		port map (
			m0_clk           => clk_clk,                                                       --   m0_clk.clk
			m0_reset         => rst_controller_reset_out_reset,                                -- m0_reset.reset
			s0_clk           => pll_100_outclk0_clk,                                           --   s0_clk.clk
			s0_reset         => rst_controller_003_reset_out_reset,                            -- s0_reset.reset
			s0_waitrequest   => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_waitrequest,   --       s0.waitrequest
			s0_readdata      => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdata,      --         .readdata
			s0_readdatavalid => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdatavalid, --         .readdatavalid
			s0_burstcount    => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_burstcount,    --         .burstcount
			s0_writedata     => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_writedata,     --         .writedata
			s0_address       => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_address,       --         .address
			s0_write         => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_write,         --         .write
			s0_read          => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_read,          --         .read
			s0_byteenable    => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_byteenable,    --         .byteenable
			s0_debugaccess   => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_debugaccess,   --         .debugaccess
			m0_waitrequest   => mm_clock_crossing_bridge_0_m0_waitrequest,                     --       m0.waitrequest
			m0_readdata      => mm_clock_crossing_bridge_0_m0_readdata,                        --         .readdata
			m0_readdatavalid => mm_clock_crossing_bridge_0_m0_readdatavalid,                   --         .readdatavalid
			m0_burstcount    => mm_clock_crossing_bridge_0_m0_burstcount,                      --         .burstcount
			m0_writedata     => mm_clock_crossing_bridge_0_m0_writedata,                       --         .writedata
			m0_address       => mm_clock_crossing_bridge_0_m0_address,                         --         .address
			m0_write         => mm_clock_crossing_bridge_0_m0_write,                           --         .write
			m0_read          => mm_clock_crossing_bridge_0_m0_read,                            --         .read
			m0_byteenable    => mm_clock_crossing_bridge_0_m0_byteenable,                      --         .byteenable
			m0_debugaccess   => mm_clock_crossing_bridge_0_m0_debugaccess                      --         .debugaccess
		);

	tightly_coupled_data_memory : component nios2_c_tightly_coupled_data_memory
		port map (
			clk        => clk_clk,                                                     --   clk1.clk
			address    => mm_interconnect_3_tightly_coupled_data_memory_s1_address,    --     s1.address
			clken      => mm_interconnect_3_tightly_coupled_data_memory_s1_clken,      --       .clken
			chipselect => mm_interconnect_3_tightly_coupled_data_memory_s1_chipselect, --       .chipselect
			write      => mm_interconnect_3_tightly_coupled_data_memory_s1_write,      --       .write
			readdata   => mm_interconnect_3_tightly_coupled_data_memory_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_3_tightly_coupled_data_memory_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_3_tightly_coupled_data_memory_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                              -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req                           --       .reset_req
		);

	key : component nios2_c_key
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_1_key_s1_address,             --                  s1.address
			write_n    => mm_interconnect_1_key_s1_write_ports_inv,     --                    .write_n
			writedata  => mm_interconnect_1_key_s1_writedata,           --                    .writedata
			chipselect => mm_interconnect_1_key_s1_chipselect,          --                    .chipselect
			readdata   => mm_interconnect_1_key_s1_readdata,            --                    .readdata
			in_port    => key_external_connection_export,               -- external_connection.export
			irq        => irq_mapper_receiver1_irq                      --                 irq.irq
		);

	timer_0 : component nios2_c_timer_0
		port map (
			clk        => clk_clk,                                      --   clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, -- reset.reset_n
			address    => mm_interconnect_1_timer_0_s1_address,         --    s1.address
			writedata  => mm_interconnect_1_timer_0_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_1_timer_0_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_1_timer_0_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_1_timer_0_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver2_irq                      --   irq.irq
		);

	ledg : component nios2_c_ledg
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_1_ledg_s1_address,            --                  s1.address
			write_n    => mm_interconnect_1_ledg_s1_write_ports_inv,    --                    .write_n
			writedata  => mm_interconnect_1_ledg_s1_writedata,          --                    .writedata
			chipselect => mm_interconnect_1_ledg_s1_chipselect,         --                    .chipselect
			readdata   => mm_interconnect_1_ledg_s1_readdata,           --                    .readdata
			out_port   => ledg_external_connection_export               -- external_connection.export
		);

	to_hex : component nios2_c_to_hex
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_1_to_hex_s1_address,          --                  s1.address
			write_n    => mm_interconnect_1_to_hex_s1_write_ports_inv,  --                    .write_n
			writedata  => mm_interconnect_1_to_hex_s1_writedata,        --                    .writedata
			chipselect => mm_interconnect_1_to_hex_s1_chipselect,       --                    .chipselect
			readdata   => mm_interconnect_1_to_hex_s1_readdata,         --                    .readdata
			out_port   => to_hex_external_connection_export             -- external_connection.export
		);

	mm_interconnect_0 : component nios2_c_mm_interconnect_0
		port map (
			clk_0_clk_clk                                                         => clk_clk,                                                            --                                                       clk_0_clk.clk
			pll_100_outclk0_clk                                                   => pll_100_outclk0_clk,                                                --                                                 pll_100_outclk0.clk
			cpu_reset_n_reset_bridge_in_reset_reset                               => rst_controller_reset_out_reset,                                     --                               cpu_reset_n_reset_bridge_in_reset.reset
			jtag_uart_reset_reset_bridge_in_reset_reset                           => rst_controller_002_reset_out_reset,                                 --                           jtag_uart_reset_reset_bridge_in_reset.reset
			mm_clock_crossing_bridge_0_s0_reset_reset_bridge_in_reset_reset       => rst_controller_003_reset_out_reset,                                 --       mm_clock_crossing_bridge_0_s0_reset_reset_bridge_in_reset.reset
			tightly_coupled_instruction_memory_reset2_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                                 -- tightly_coupled_instruction_memory_reset2_reset_bridge_in_reset.reset
			cpu_data_master_address                                               => cpu_data_master_address,                                            --                                                 cpu_data_master.address
			cpu_data_master_waitrequest                                           => cpu_data_master_waitrequest,                                        --                                                                .waitrequest
			cpu_data_master_burstcount                                            => cpu_data_master_burstcount,                                         --                                                                .burstcount
			cpu_data_master_byteenable                                            => cpu_data_master_byteenable,                                         --                                                                .byteenable
			cpu_data_master_read                                                  => cpu_data_master_read,                                               --                                                                .read
			cpu_data_master_readdata                                              => cpu_data_master_readdata,                                           --                                                                .readdata
			cpu_data_master_readdatavalid                                         => cpu_data_master_readdatavalid,                                      --                                                                .readdatavalid
			cpu_data_master_write                                                 => cpu_data_master_write,                                              --                                                                .write
			cpu_data_master_writedata                                             => cpu_data_master_writedata,                                          --                                                                .writedata
			cpu_data_master_debugaccess                                           => cpu_data_master_debugaccess,                                        --                                                                .debugaccess
			cpu_instruction_master_address                                        => cpu_instruction_master_address,                                     --                                          cpu_instruction_master.address
			cpu_instruction_master_waitrequest                                    => cpu_instruction_master_waitrequest,                                 --                                                                .waitrequest
			cpu_instruction_master_burstcount                                     => cpu_instruction_master_burstcount,                                  --                                                                .burstcount
			cpu_instruction_master_read                                           => cpu_instruction_master_read,                                        --                                                                .read
			cpu_instruction_master_readdata                                       => cpu_instruction_master_readdata,                                    --                                                                .readdata
			cpu_instruction_master_readdatavalid                                  => cpu_instruction_master_readdatavalid,                               --                                                                .readdatavalid
			cpu_jtag_debug_module_address                                         => mm_interconnect_0_cpu_jtag_debug_module_address,                    --                                           cpu_jtag_debug_module.address
			cpu_jtag_debug_module_write                                           => mm_interconnect_0_cpu_jtag_debug_module_write,                      --                                                                .write
			cpu_jtag_debug_module_read                                            => mm_interconnect_0_cpu_jtag_debug_module_read,                       --                                                                .read
			cpu_jtag_debug_module_readdata                                        => mm_interconnect_0_cpu_jtag_debug_module_readdata,                   --                                                                .readdata
			cpu_jtag_debug_module_writedata                                       => mm_interconnect_0_cpu_jtag_debug_module_writedata,                  --                                                                .writedata
			cpu_jtag_debug_module_byteenable                                      => mm_interconnect_0_cpu_jtag_debug_module_byteenable,                 --                                                                .byteenable
			cpu_jtag_debug_module_waitrequest                                     => mm_interconnect_0_cpu_jtag_debug_module_waitrequest,                --                                                                .waitrequest
			cpu_jtag_debug_module_debugaccess                                     => mm_interconnect_0_cpu_jtag_debug_module_debugaccess,                --                                                                .debugaccess
			jtag_uart_avalon_jtag_slave_address                                   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,              --                                     jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write                                     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,                --                                                                .write
			jtag_uart_avalon_jtag_slave_read                                      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,                 --                                                                .read
			jtag_uart_avalon_jtag_slave_readdata                                  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,             --                                                                .readdata
			jtag_uart_avalon_jtag_slave_writedata                                 => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,            --                                                                .writedata
			jtag_uart_avalon_jtag_slave_waitrequest                               => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,          --                                                                .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                                => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,           --                                                                .chipselect
			mm_clock_crossing_bridge_0_s0_address                                 => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_address,            --                                   mm_clock_crossing_bridge_0_s0.address
			mm_clock_crossing_bridge_0_s0_write                                   => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_write,              --                                                                .write
			mm_clock_crossing_bridge_0_s0_read                                    => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_read,               --                                                                .read
			mm_clock_crossing_bridge_0_s0_readdata                                => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdata,           --                                                                .readdata
			mm_clock_crossing_bridge_0_s0_writedata                               => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_writedata,          --                                                                .writedata
			mm_clock_crossing_bridge_0_s0_burstcount                              => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_burstcount,         --                                                                .burstcount
			mm_clock_crossing_bridge_0_s0_byteenable                              => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_byteenable,         --                                                                .byteenable
			mm_clock_crossing_bridge_0_s0_readdatavalid                           => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdatavalid,      --                                                                .readdatavalid
			mm_clock_crossing_bridge_0_s0_waitrequest                             => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_waitrequest,        --                                                                .waitrequest
			mm_clock_crossing_bridge_0_s0_debugaccess                             => mm_interconnect_0_mm_clock_crossing_bridge_0_s0_debugaccess,        --                                                                .debugaccess
			sysid_qsys_0_control_slave_address                                    => mm_interconnect_0_sysid_qsys_0_control_slave_address,               --                                      sysid_qsys_0_control_slave.address
			sysid_qsys_0_control_slave_readdata                                   => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,              --                                                                .readdata
			tightly_coupled_instruction_memory_s2_address                         => mm_interconnect_0_tightly_coupled_instruction_memory_s2_address,    --                           tightly_coupled_instruction_memory_s2.address
			tightly_coupled_instruction_memory_s2_write                           => mm_interconnect_0_tightly_coupled_instruction_memory_s2_write,      --                                                                .write
			tightly_coupled_instruction_memory_s2_readdata                        => mm_interconnect_0_tightly_coupled_instruction_memory_s2_readdata,   --                                                                .readdata
			tightly_coupled_instruction_memory_s2_writedata                       => mm_interconnect_0_tightly_coupled_instruction_memory_s2_writedata,  --                                                                .writedata
			tightly_coupled_instruction_memory_s2_byteenable                      => mm_interconnect_0_tightly_coupled_instruction_memory_s2_byteenable, --                                                                .byteenable
			tightly_coupled_instruction_memory_s2_chipselect                      => mm_interconnect_0_tightly_coupled_instruction_memory_s2_chipselect, --                                                                .chipselect
			tightly_coupled_instruction_memory_s2_clken                           => mm_interconnect_0_tightly_coupled_instruction_memory_s2_clken       --                                                                .clken
		);

	mm_interconnect_1 : component nios2_c_mm_interconnect_1
		port map (
			clk_0_clk_clk                                                   => clk_clk,                                     --                                                 clk_0_clk.clk
			key_reset_reset_bridge_in_reset_reset                           => rst_controller_001_reset_out_reset,          --                           key_reset_reset_bridge_in_reset.reset
			mm_clock_crossing_bridge_0_m0_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,              -- mm_clock_crossing_bridge_0_m0_reset_reset_bridge_in_reset.reset
			mm_clock_crossing_bridge_0_m0_address                           => mm_clock_crossing_bridge_0_m0_address,       --                             mm_clock_crossing_bridge_0_m0.address
			mm_clock_crossing_bridge_0_m0_waitrequest                       => mm_clock_crossing_bridge_0_m0_waitrequest,   --                                                          .waitrequest
			mm_clock_crossing_bridge_0_m0_burstcount                        => mm_clock_crossing_bridge_0_m0_burstcount,    --                                                          .burstcount
			mm_clock_crossing_bridge_0_m0_byteenable                        => mm_clock_crossing_bridge_0_m0_byteenable,    --                                                          .byteenable
			mm_clock_crossing_bridge_0_m0_read                              => mm_clock_crossing_bridge_0_m0_read,          --                                                          .read
			mm_clock_crossing_bridge_0_m0_readdata                          => mm_clock_crossing_bridge_0_m0_readdata,      --                                                          .readdata
			mm_clock_crossing_bridge_0_m0_readdatavalid                     => mm_clock_crossing_bridge_0_m0_readdatavalid, --                                                          .readdatavalid
			mm_clock_crossing_bridge_0_m0_write                             => mm_clock_crossing_bridge_0_m0_write,         --                                                          .write
			mm_clock_crossing_bridge_0_m0_writedata                         => mm_clock_crossing_bridge_0_m0_writedata,     --                                                          .writedata
			mm_clock_crossing_bridge_0_m0_debugaccess                       => mm_clock_crossing_bridge_0_m0_debugaccess,   --                                                          .debugaccess
			key_s1_address                                                  => mm_interconnect_1_key_s1_address,            --                                                    key_s1.address
			key_s1_write                                                    => mm_interconnect_1_key_s1_write,              --                                                          .write
			key_s1_readdata                                                 => mm_interconnect_1_key_s1_readdata,           --                                                          .readdata
			key_s1_writedata                                                => mm_interconnect_1_key_s1_writedata,          --                                                          .writedata
			key_s1_chipselect                                               => mm_interconnect_1_key_s1_chipselect,         --                                                          .chipselect
			ledg_s1_address                                                 => mm_interconnect_1_ledg_s1_address,           --                                                   ledg_s1.address
			ledg_s1_write                                                   => mm_interconnect_1_ledg_s1_write,             --                                                          .write
			ledg_s1_readdata                                                => mm_interconnect_1_ledg_s1_readdata,          --                                                          .readdata
			ledg_s1_writedata                                               => mm_interconnect_1_ledg_s1_writedata,         --                                                          .writedata
			ledg_s1_chipselect                                              => mm_interconnect_1_ledg_s1_chipselect,        --                                                          .chipselect
			timer_0_s1_address                                              => mm_interconnect_1_timer_0_s1_address,        --                                                timer_0_s1.address
			timer_0_s1_write                                                => mm_interconnect_1_timer_0_s1_write,          --                                                          .write
			timer_0_s1_readdata                                             => mm_interconnect_1_timer_0_s1_readdata,       --                                                          .readdata
			timer_0_s1_writedata                                            => mm_interconnect_1_timer_0_s1_writedata,      --                                                          .writedata
			timer_0_s1_chipselect                                           => mm_interconnect_1_timer_0_s1_chipselect,     --                                                          .chipselect
			to_hex_s1_address                                               => mm_interconnect_1_to_hex_s1_address,         --                                                 to_hex_s1.address
			to_hex_s1_write                                                 => mm_interconnect_1_to_hex_s1_write,           --                                                          .write
			to_hex_s1_readdata                                              => mm_interconnect_1_to_hex_s1_readdata,        --                                                          .readdata
			to_hex_s1_writedata                                             => mm_interconnect_1_to_hex_s1_writedata,       --                                                          .writedata
			to_hex_s1_chipselect                                            => mm_interconnect_1_to_hex_s1_chipselect       --                                                          .chipselect
		);

	mm_interconnect_2 : component nios2_c_mm_interconnect_2
		port map (
			clk_0_clk_clk                                          => clk_clk,                                                            --                                clk_0_clk.clk
			cpu_reset_n_reset_bridge_in_reset_reset                => rst_controller_reset_out_reset,                                     --        cpu_reset_n_reset_bridge_in_reset.reset
			cpu_tightly_coupled_instruction_master_0_address       => cpu_tightly_coupled_instruction_master_0_address,                   -- cpu_tightly_coupled_instruction_master_0.address
			cpu_tightly_coupled_instruction_master_0_waitrequest   => cpu_tightly_coupled_instruction_master_0_waitrequest,               --                                         .waitrequest
			cpu_tightly_coupled_instruction_master_0_read          => cpu_tightly_coupled_instruction_master_0_read,                      --                                         .read
			cpu_tightly_coupled_instruction_master_0_readdata      => cpu_tightly_coupled_instruction_master_0_readdata,                  --                                         .readdata
			cpu_tightly_coupled_instruction_master_0_readdatavalid => cpu_tightly_coupled_instruction_master_0_readdatavalid,             --                                         .readdatavalid
			cpu_tightly_coupled_instruction_master_0_clken         => cpu_tightly_coupled_instruction_master_0_clken,                     --                                         .clken
			tightly_coupled_instruction_memory_s1_address          => mm_interconnect_2_tightly_coupled_instruction_memory_s1_address,    --    tightly_coupled_instruction_memory_s1.address
			tightly_coupled_instruction_memory_s1_write            => mm_interconnect_2_tightly_coupled_instruction_memory_s1_write,      --                                         .write
			tightly_coupled_instruction_memory_s1_readdata         => mm_interconnect_2_tightly_coupled_instruction_memory_s1_readdata,   --                                         .readdata
			tightly_coupled_instruction_memory_s1_writedata        => mm_interconnect_2_tightly_coupled_instruction_memory_s1_writedata,  --                                         .writedata
			tightly_coupled_instruction_memory_s1_byteenable       => mm_interconnect_2_tightly_coupled_instruction_memory_s1_byteenable, --                                         .byteenable
			tightly_coupled_instruction_memory_s1_chipselect       => mm_interconnect_2_tightly_coupled_instruction_memory_s1_chipselect, --                                         .chipselect
			tightly_coupled_instruction_memory_s1_clken            => mm_interconnect_2_tightly_coupled_instruction_memory_s1_clken       --                                         .clken
		);

	mm_interconnect_3 : component nios2_c_mm_interconnect_3
		port map (
			clk_0_clk_clk                                   => clk_clk,                                                     --                         clk_0_clk.clk
			cpu_reset_n_reset_bridge_in_reset_reset         => rst_controller_reset_out_reset,                              -- cpu_reset_n_reset_bridge_in_reset.reset
			cpu_tightly_coupled_data_master_0_address       => cpu_tightly_coupled_data_master_0_address,                   -- cpu_tightly_coupled_data_master_0.address
			cpu_tightly_coupled_data_master_0_waitrequest   => cpu_tightly_coupled_data_master_0_waitrequest,               --                                  .waitrequest
			cpu_tightly_coupled_data_master_0_byteenable    => cpu_tightly_coupled_data_master_0_byteenable,                --                                  .byteenable
			cpu_tightly_coupled_data_master_0_read          => cpu_tightly_coupled_data_master_0_read,                      --                                  .read
			cpu_tightly_coupled_data_master_0_readdata      => cpu_tightly_coupled_data_master_0_readdata,                  --                                  .readdata
			cpu_tightly_coupled_data_master_0_readdatavalid => cpu_tightly_coupled_data_master_0_readdatavalid,             --                                  .readdatavalid
			cpu_tightly_coupled_data_master_0_write         => cpu_tightly_coupled_data_master_0_write,                     --                                  .write
			cpu_tightly_coupled_data_master_0_writedata     => cpu_tightly_coupled_data_master_0_writedata,                 --                                  .writedata
			cpu_tightly_coupled_data_master_0_clken         => cpu_tightly_coupled_data_master_0_clken,                     --                                  .clken
			tightly_coupled_data_memory_s1_address          => mm_interconnect_3_tightly_coupled_data_memory_s1_address,    --    tightly_coupled_data_memory_s1.address
			tightly_coupled_data_memory_s1_write            => mm_interconnect_3_tightly_coupled_data_memory_s1_write,      --                                  .write
			tightly_coupled_data_memory_s1_readdata         => mm_interconnect_3_tightly_coupled_data_memory_s1_readdata,   --                                  .readdata
			tightly_coupled_data_memory_s1_writedata        => mm_interconnect_3_tightly_coupled_data_memory_s1_writedata,  --                                  .writedata
			tightly_coupled_data_memory_s1_byteenable       => mm_interconnect_3_tightly_coupled_data_memory_s1_byteenable, --                                  .byteenable
			tightly_coupled_data_memory_s1_chipselect       => mm_interconnect_3_tightly_coupled_data_memory_s1_chipselect, --                                  .chipselect
			tightly_coupled_data_memory_s1_clken            => mm_interconnect_3_tightly_coupled_data_memory_s1_clken       --                                  .clken
		);

	irq_mapper : component nios2_c_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			sender_irq    => cpu_d_irq_irq                   --    sender.irq
		);

	irq_synchronizer : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => pll_100_outclk0_clk,                --       receiver_clk.clk
			sender_clk     => clk_clk,                            --         sender_clk.clk
			receiver_reset => rst_controller_002_reset_out_reset, -- receiver_clk_reset.reset
			sender_reset   => rst_controller_reset_out_reset,     --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_receiver_irq,      --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver0_irq            --             sender.irq
		);

	rst_controller : component nios2_c_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => cpu_jtag_debug_module_reset_reset,  -- reset_in1.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_001 : component nios2_c_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			clk            => clk_clk,                                --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_001_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_in1      => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_002 : component nios2_c_rst_controller_002
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => cpu_jtag_debug_module_reset_reset,  -- reset_in1.reset
			clk            => pll_100_outclk0_clk,                --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_003 : component nios2_c_rst_controller_003
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => pll_100_outclk0_clk,                --       clk.clk
			reset_out      => rst_controller_003_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_1_to_hex_s1_write_ports_inv <= not mm_interconnect_1_to_hex_s1_write;

	mm_interconnect_1_key_s1_write_ports_inv <= not mm_interconnect_1_key_s1_write;

	mm_interconnect_1_ledg_s1_write_ports_inv <= not mm_interconnect_1_ledg_s1_write;

	mm_interconnect_1_timer_0_s1_write_ports_inv <= not mm_interconnect_1_timer_0_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

	rst_controller_002_reset_out_reset_ports_inv <= not rst_controller_002_reset_out_reset;

end architecture rtl; -- of nios2_c
